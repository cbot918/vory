module main

import vory

fn main() {
	v := vory.new_vory()
	v.hello()
}
