module model

pub struct Users{
pub mut:
	id string
	name string
	email string
}